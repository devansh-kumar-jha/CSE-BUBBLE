`include "../../source/processor.v"

module bubble_sort_test();
    // Program in form of Instructions loaded into the Instruction Memory

    // Instantiate the Processor Module

    // Upon getting signal from processor finish the simulation
    // call $finish;

endmodule
