/// This will be a combinational logic.
module transfer(initial_pc,r0,r1,const,pc);
    input [31:0] initial_pc,r0,r1,const;
    output [31:0] pc;

    // reg [31:0] pc_check;
    // wire [4:0] r0,r1,r2;
    // assign r1 = ir[25:21];
    // assign r0 = ir[20:16];
    // assign num = ir[15:0];

    // always @(*) begin
    //     check <= data_in;
    // end

    // assign data_out <= check;
endmodule