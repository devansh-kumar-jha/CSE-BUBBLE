//! These are the memory modules which will be called and used in the processor module. They all will be present in the
//! write mode until the loading phase of the processor is running after that instruction memory would convert into
//! read only mode but the data memory would still be present in write mode to the user.

/// This is the module which will be used as the source of memory and this has the following controls as explained
// clk - The synchronizing signal for all the phases of the processor machine.
// reset - The reset signal to delete and restart the whole memory.
// in - The data which is send as input for storing in memory.
// out - The data which is being asked for from memory.
// mode - The working mode of the memory currently. 0 means write mode and 1 means read only mode.
// address_a - The address at which the input is filled by the memory.
// address_b - The address from which output is generated by the memory.
// writeEnable - In write mode when we have to refrain from writing into memory disable this flag.
module veda_instruction #(parameter width = 32, parameter depth = 256, parameter len = 8) (clk,reset,in,out,mode,address_a,address_b,writeEnable);
    input wire [width-1:0] in;
    input wire [len-1:0] address_a,address_b;
    input wire clk,reset,mode,writeEnable;                                // Mode 0 means write mode and Mode 1 means read mode
    output wire [width-1:0] out;
    
    reg [width-1:0] memory[0:depth-1];
    reg [width-1:0] dataout,cur;
    integer i;

    // Setting the memory at erased state.
    initial begin
        cur <= 0;
    end

    initial begin
        #1
        // Write program to enter instruction memory into the machine
        memory[0]  <= 32'b001000_00110_11011_0000000000000000;               // lw $27, 0($6)  $s3 = 10
        memory[0]  <= 32'b000001_00110_11010_0000000000000001;               // addi $26, $6, 1  $s2 = 1
        memory[0]  <= 32'b000000_00110_10001_0000000000000000;               // addi $17, $6, 0
        memory[1]  <= 32'b000000_11011_10001_10010_00000_000001;             // sub $18, $27, $17
        memory[2]  <= 32'b000001_10010_10010_1111111111111111;               // addi $18, $18, -1
        memory[3]  <= 32'b000001_00110_10011_0000000000000000;               // addi $19, $6, 0
        memory[4]  <= 32'b000000_10011_10010_11001_00000_000001;             // sub $25, $19, $18
        memory[5]  <= 32'b010011_11001_00110_11111_00000_000000;             // slt $31, $25, $6
        memory[6]  <= 32'b001010_00110_11111_0000000000001101;               // beq $31, $6, 13
        memory[7]  <= 32'b001101_00110_11001_0000000000001100;               // bgte $25, $6, 12
        memory[8]  <= 32'b000111_10011_10100_0000000000000010;               // sll $20, $19, 2
        memory[9]  <= 32'b000000_10100_11000_10100_00000_000000;
        memory[10] <= 32'b000000_10100_10101_0000000000000100;
        memory[11] <= 32'b001000_10100_10110_0000000000000000;
        memory[12] <= 32'b001000_10101_10111_0000000000000000;
        memory[13] <= 32'b000000_10110_10111_11000_00000_000001;
        memory[14] <= 32'b010011_11000_00110_11111_00000_000000;
        memory[15] <= 32'b001011_00110_11111_0000000000000011;
        memory[16] <= 32'b001001_10101_10110_0000000000000000;
        memory[17] <= 32'b001001_10100_10111_0000000000000000;
        memory[18] <= 32'b000000_10011_10011_0000000000000001;
        memory[19] <= 32'b001011_10010_10011_1111111111110101;   
        memory[20] <= 32'b000000_10001_10001_0000000000000001;
        memory[21] <= 32'b001011_11001_10011_1111111111101100;
        memory[22] <= 32'b100001_00000000000000000000010000;
        cur <= 23;
    end
    
    // Sequential write operation at posedge of clk.
    always @(posedge reset or posedge clk) begin
        if(reset==1'b1) begin
            dataout <= 0;
            for(i=cur;i<depth;i=i+1) begin memory[i] <= 0; end
        end
        else begin
            if(writeEnable==1'b1 && mode==1'b0) begin
                memory[address_a] <= in;
            end
        end
    end

    // Combinational read operation.
    assign out = memory[address_b];
endmodule


/// This is the module which will be used as the source of memory and this has the following controls as explained
// clk - The synchronizing signal for all the phases of the processor machine.
// reset - The reset signal to delete and restart the whole memory.
// in - The data which is send as input for storing in memory.
// out - The data which is being asked for from memory.
// mode - The working mode of the memory currently. 0 means write mode and 1 means read only mode.
// address_a - The address at which the input is filled by the memory.
// address_b - The address from which output is generated by the memory.
// writeEnable - In write mode when we have to refrain from writing into memory disable this flag.
module veda_data #(parameter width = 32, parameter depth = 256, parameter len = 8) (clk,reset,in,out,mode,address_a,address_b,writeEnable);
    input wire [width-1:0] in;
    input wire [len-1:0] address_a,address_b;
    input wire clk,reset,mode,writeEnable;                            // Mode 0 means write mode and Mode 1 means read mode
    output wire [width-1:0] out;
    
    reg [width-1:0] memory[0:depth-1];
    reg [width-1:0] dataout,cur;
    integer i;

    // Setting the memory at erased state.
    initial begin
        cur <= 0;
    end
    
    initial begin
        #1
        // Write program to enter data memory into the machine
        memory[0] <= 32'd10;                        // Length of array
        memory[1] <= 32'd643;                       // Starting address of array in data memory
        memory[2] <= 32'd573;
        memory[3] <= 32'd532;
        memory[4] <= 32'd087;
        memory[5] <= 32'd879;
        memory[6] <= 32'd242;
        memory[7] <= 32'd64;
        memory[8] <= 32'd805;
        memory[9] <= 32'd868;
        memory[10] <= 32'd57320;
        memory[11] <= 32'd378;                      // Last value in array to be sorted
        cur <= 12;
    end
    
    // Sequential write operation at posedge of clk.
    always @(posedge reset or posedge clk) begin
        if(reset==1'b1) begin
            dataout <= 0;
            for(i=cur;i<depth;i=i+1) begin memory[i] <= 0; end
        end
        else begin
            if(writeEnable==1'b1 && mode==1'b0) begin
                memory[address_a] <= in;
            end
        end
    end

    // Combinational read operation.
    assign out = memory[address_b];
endmodule
