// This file will run the Instruction Fetch phase inside the processor.
// Here in the instruction will be loaded inside the Instruction Register in 1 clock cycle
// The module takes input the program counter and the instruction memory from the processor
// and outputs the instruction in IR register

module instr_fetch();

endmodule
