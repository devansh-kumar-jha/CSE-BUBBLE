//! These are the memory modules which will be called and used in the processor module. They all will be present in the
//! write mode until the loading phase of the processor is running after that instruction memory would convert into
//! read only mode but the data memory would still be present in write mode to the user.

/// This is the module which will be used as the source of memory and this has the following controls as explained
// clk - The synchronizing signal for all the phases of the processor machine.
// reset - The reset signal to delete and restart the whole memory.
// in - The data which is send as input for storing in memory.
// out - The data which is being asked for from memory.
// mode - The working mode of the memory currently. 0 means write mode and 1 means read only mode.
// address_a - The address at which the input is filled by the memory.
// address_b - The address from which output is generated by the memory.
// writeEnable - In write mode when we have to refrain from writing into memory disable this flag.
module veda #(parameter width = 32, parameter depth = 256, parameter len = 8) (clk,reset,in,out,mode,address_a,address_b,writeEnable);
    input wire [width-1:0] in;
    input wire [len-1:0] address_a,address_b;
    input wire clk,reset,mode,writeEnable; // Mode 0 means write mode and Mode 1 means read mode
    output wire [width-1:0] out;
    
    reg [width-1:0] memory[0:depth-1];
    reg [width-1:0] dataout;
    integer i;

    // initial begin
    //     memory[0] <= 32'b000001_00110_10101_0000000011111111;                      // addi $t4, $0, num1
    //     memory[1] <= 32'b000001_00110_10110_0000000011111110;                      // addi $t5, $0, num2
    //     memory[2] <= 32'b000001_00110_10111_0000000011111101;                      // addi $t6, $0, num3
    //     memory[3] <= 32'b001000_10101_10001_0000000000000000;                      // lw $t0, 0($t4)
    //     memory[4] <= 32'b001000_10110_10010_0000000000000000;                      // lw $t1, 0($t5)
    //     memory[5] <= 32'b001000_10111_10011_0000000000000000;                      // lw $t2, 0($t6)
    //     memory[6] <= 32'b000000_10011_10010_10101_00000_000001;                    // sub $t4, $t2, $t1
    //     memory[7] <= 32'b000001_00110_01000_0000000000000001;                      // loopp1: addi $v0, $0, 1
    //     memory[8] <= 32'b000001_10101_01010_0000000000000000;                      // addi $a0, $t4, 0
    //     memory[9] <= 32'b010101_00000000000000000000000000;                        // syscall
    //     memory[10] <= 32'b000001_10101_10101_0000000000000001;                     // addi $t4, $t4, 1
    //     // #10 new_instruction <= 32'b001000_00010_00001_0000000000001100;         // bne $t4, $t0, loopp1
    //     memory[11] <= 32'b000001_00110_01000_0000000000000010;                     // addi $v0, $0, 2
    //     memory[12] <= 32'b010101_00000000000000000000000000;                       // syscall
    // end
    
    // Sequential write operation at posedge of clk.
    always @(posedge reset or posedge clk) begin
        if(reset==1'b1) begin
            dataout <= 0;
            for(i=0;i<depth;i=i+1) begin memory[i] <= 0; end
        end
        else begin
            if(writeEnable==1'b1 && mode==1'b0) begin
                memory[address_a] <= in;
            end
        end
    end

    // Combinational read operation.
    assign out = memory[address_b];
endmodule

/// This is the module which will be used as the source of memory and this has the following controls as explained
// clk - The synchronizing signal for all the phases of the processor machine.
// reset - The reset signal to delete and restart the whole memory.
// in - The data which is send as input for storing in memory.
// out - The data which is being asked for from memory.
// mode - The working mode of the memory currently. 0 means write mode and 1 means read only mode.
// address_a - The address at which the input is filled by the memory.
// address_b - The address from which output is generated by the memory.
// writeEnable - In write mode when we have to refrain from writing into memory disable this flag.
module veda_data #(parameter width = 32, parameter depth = 256, parameter len = 8) (clk,reset,in,out,mode,address_a,address_b,writeEnable);
    input wire [width-1:0] in;
    input wire [len-1:0] address_a,address_b;
    input wire clk,reset,mode,writeEnable; // Mode 0 means write mode and Mode 1 means read mode
    output wire [width-1:0] out;
    
    reg [width-1:0] memory[0:depth-1];
    reg [width-1:0] dataout;
    integer i;

    // initial begin
    //     memory[0] <= 32'b00000000000000000000000000001010;                     // num1:   .word 10 stored at data[255]
    //     memory[1] <= 32'b00000000000000000000000000000110;                     // num2:   .word 6 stored at data[254]
    //     memory[2] <= 32'b00000000000000000000000000001101;                     // num3:   .word 13 stored at data[253]
    // end
    
    // Sequential write operation at posedge of clk.
    always @(posedge reset or posedge clk) begin
        if(reset==1'b1) begin
            dataout <= 0;
            for(i=0;i<depth;i=i+1) begin memory[i] <= 0; end
        end
        else begin
            if(writeEnable==1'b1 && mode==1'b0) begin
                memory[address_a] <= in;
            end
        end
    end

    // Combinational read operation.
    assign out = memory[address_b];
endmodule
