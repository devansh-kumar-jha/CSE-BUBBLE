//! These are the memory modules which will be called and used in the processor module. They all will be present in the
//! write mode until the loading phase of the processor is running after that instruction memory would convert into
//! read only mode but the data memory would still be present in write mode to the user.

/// This is the module which will be used as the source of memory and this has the following controls as explained
// clk - The synchronizing signal for all the phases of the processor machine.
// reset - The reset signal to delete and restart the whole memory.
// in - The data which is send as input for storing in memory.
// out - The data which is being asked for from memory.
// mode - The working mode of the memory currently. 0 means write mode and 1 means read only mode.
// address_a - The address at which the input is filled by the memory.
// address_b - The address from which output is generated by the memory.
// writeEnable - In write mode when we have to refrain from writing into memory disable this flag.
module veda #(parameter width = 32, parameter depth = 256, parameter len = 8) (clk,reset,in,out,mode,address_a,address_b,writeEnable);
    input wire [width-1:0] in;
    input wire [len-1:0] address_a,address_b;
    input wire clk,reset,mode,writeEnable; // Mode 0 means write mode and Mode 1 means read mode
    output wire [width-1:0] out;
    
    reg [width-1:0] memory[0:depth-1];
    reg [width-1:0] dataout;
    integer i;

    always @(posedge reset or posedge clk) begin
        if(reset==1'b1) begin
            dataout <= 0;
            for(i=0;i<depth;i=i+1) begin memory[i] <= 0; end
        end
        else begin
            if(writeEnable==1'b1 && mode==1'b0) begin
                memory[address_a] = in;
            end
            dataout = memory[address_b];
        end
    end
    assign out = dataout;
endmodule
